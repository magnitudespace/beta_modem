module filter8(
  input CLK,
  input ENABLE,
  input [3:0] STAGE,//should be parametrized size 
  input [65:0] INPUT_I,//should be parametrized size 
  input [65:0] INPUT_Q,//should be parametrized size 
  output [12:0] OUTPUT_I,
  output [12:0] OUTPUT_Q
);

  wire [13:0] sum;
  reg signed [12:0] result_i = 0;
  reg signed [12:0] result_q = 0;

  assign OUTPUT_I = result_i;
  assign OUTPUT_Q = result_q;

  wire [65:0] INPUT;//should be parametrized size 

  assign INPUT = STAGE[0] ? INPUT_Q : INPUT_I;

reg [13:0] a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a20, a21, a22, a23, a24, a25, a26, a27, a28, a29, a30, a31, a32;

always @ (STAGE or INPUT) 
begin

  a0 = 0;
  case ({STAGE[3:1], INPUT[1:0]})
    5'b00000 : a0 = 0;
    5'b00001 : a0 = -3;
    5'b00010 : a0 = 0;
    5'b00011 : a0 = 3;
    5'b00100 : a0 = 0;
    5'b00101 : a0 = 0;
    5'b00110 : a0 = 0;
    5'b00111 : a0 = 0;
    5'b01000 : a0 = 0;
    5'b01001 : a0 = 0;
    5'b01010 : a0 = 0;
    5'b01011 : a0 = 0;
    5'b01100 : a0 = 0;
    5'b01101 : a0 = 0;
    5'b01110 : a0 = 0;
    5'b01111 : a0 = 0;
    5'b10000 : a0 = 0;
    5'b10001 : a0 = 0;
    5'b10010 : a0 = 0;
    5'b10011 : a0 = 0;
    5'b10100 : a0 = 0;
    5'b10101 : a0 = 0;
    5'b10110 : a0 = 0;
    5'b10111 : a0 = 0;
    5'b11000 : a0 = 0;
    5'b11001 : a0 = 0;
    5'b11010 : a0 = 0;
    5'b11011 : a0 = 0;
    5'b11100 : a0 = 0;
    5'b11101 : a0 = 0;
    5'b11110 : a0 = 0;
    5'b11111 : a0 = 0;
  endcase

  a1 = 0;
  case ({STAGE[3:1], INPUT[3:2]})
    5'b00000 : a1 = 0;
    5'b00001 : a1 = 0;
    5'b00010 : a1 = 0;
    5'b00011 : a1 = 0;
    5'b00100 : a1 = 0;
    5'b00101 : a1 = 2;
    5'b00110 : a1 = 0;
    5'b00111 : a1 = -2;
    5'b01000 : a1 = 0;
    5'b01001 : a1 = 5;
    5'b01010 : a1 = 0;
    5'b01011 : a1 = -5;
    5'b01100 : a1 = 0;
    5'b01101 : a1 = 6;
    5'b01110 : a1 = 0;
    5'b01111 : a1 = -6;
    5'b10000 : a1 = 0;
    5'b10001 : a1 = 6;
    5'b10010 : a1 = 0;
    5'b10011 : a1 = -6;
    5'b10100 : a1 = 0;
    5'b10101 : a1 = 4;
    5'b10110 : a1 = 0;
    5'b10111 : a1 = -4;
    5'b11000 : a1 = 0;
    5'b11001 : a1 = 2;
    5'b11010 : a1 = 0;
    5'b11011 : a1 = -2;
    5'b11100 : a1 = 0;
    5'b11101 : a1 = 0;
    5'b11110 : a1 = 0;
    5'b11111 : a1 = 0;
  endcase

  a2 = 0;
  case ({STAGE[3:1], INPUT[5:4]})
    5'b00000 : a2 = 0;
    5'b00001 : a2 = 5;
    5'b00010 : a2 = 0;
    5'b00011 : a2 = -5;
    5'b00100 : a2 = 0;
    5'b00101 : a2 = 2;
    5'b00110 : a2 = 0;
    5'b00111 : a2 = -2;
    5'b01000 : a2 = 0;
    5'b01001 : a2 = 0;
    5'b01010 : a2 = 0;
    5'b01011 : a2 = 0;
    5'b01100 : a2 = 0;
    5'b01101 : a2 = -3;
    5'b01110 : a2 = 0;
    5'b01111 : a2 = 3;
    5'b10000 : a2 = 0;
    5'b10001 : a2 = -6;
    5'b10010 : a2 = 0;
    5'b10011 : a2 = 6;
    5'b10100 : a2 = 0;
    5'b10101 : a2 = -6;
    5'b10110 : a2 = 0;
    5'b10111 : a2 = 6;
    5'b11000 : a2 = 0;
    5'b11001 : a2 = -5;
    5'b11010 : a2 = 0;
    5'b11011 : a2 = 5;
    5'b11100 : a2 = 0;
    5'b11101 : a2 = -3;
    5'b11110 : a2 = 0;
    5'b11111 : a2 = 3;
  endcase

  a3 = 0;
  case ({STAGE[3:1], INPUT[7:6]})
    5'b00000 : a3 = 0;
    5'b00001 : a3 = -9;
    5'b00010 : a3 = 0;
    5'b00011 : a3 = 9;
    5'b00100 : a3 = 0;
    5'b00101 : a3 = -8;
    5'b00110 : a3 = 0;
    5'b00111 : a3 = 8;
    5'b01000 : a3 = 0;
    5'b01001 : a3 = -5;
    5'b01010 : a3 = 0;
    5'b01011 : a3 = 5;
    5'b01100 : a3 = 0;
    5'b01101 : a3 = -1;
    5'b01110 : a3 = 0;
    5'b01111 : a3 = 1;
    5'b10000 : a3 = 0;
    5'b10001 : a3 = 2;
    5'b10010 : a3 = 0;
    5'b10011 : a3 = -2;
    5'b10100 : a3 = 0;
    5'b10101 : a3 = 5;
    5'b10110 : a3 = 0;
    5'b10111 : a3 = -5;
    5'b11000 : a3 = 0;
    5'b11001 : a3 = 7;
    5'b11010 : a3 = 0;
    5'b11011 : a3 = -7;
    5'b11100 : a3 = 0;
    5'b11101 : a3 = 7;
    5'b11110 : a3 = 0;
    5'b11111 : a3 = -7;
  endcase

  a4 = 0;
  case ({STAGE[3:1], INPUT[9:8]})
    5'b00000 : a4 = 0;
    5'b00001 : a4 = 8;
    5'b00010 : a4 = 0;
    5'b00011 : a4 = -8;
    5'b00100 : a4 = 0;
    5'b00101 : a4 = 10;
    5'b00110 : a4 = 0;
    5'b00111 : a4 = -10;
    5'b01000 : a4 = 0;
    5'b01001 : a4 = 10;
    5'b01010 : a4 = 0;
    5'b01011 : a4 = -10;
    5'b01100 : a4 = 0;
    5'b01101 : a4 = 8;
    5'b01110 : a4 = 0;
    5'b01111 : a4 = -8;
    5'b10000 : a4 = 0;
    5'b10001 : a4 = 4;
    5'b10010 : a4 = 0;
    5'b10011 : a4 = -4;
    5'b10100 : a4 = 0;
    5'b10101 : a4 = 0;
    5'b10110 : a4 = 0;
    5'b10111 : a4 = 0;
    5'b11000 : a4 = 0;
    5'b11001 : a4 = -4;
    5'b11010 : a4 = 0;
    5'b11011 : a4 = 4;
    5'b11100 : a4 = 0;
    5'b11101 : a4 = -7;
    5'b11110 : a4 = 0;
    5'b11111 : a4 = 7;
  endcase

  a5 = 0;
  case ({STAGE[3:1], INPUT[11:10]})
    5'b00000 : a5 = 0;
    5'b00001 : a5 = -2;
    5'b00010 : a5 = 0;
    5'b00011 : a5 = 2;
    5'b00100 : a5 = 0;
    5'b00101 : a5 = -7;
    5'b00110 : a5 = 0;
    5'b00111 : a5 = 7;
    5'b01000 : a5 = 0;
    5'b01001 : a5 = -11;
    5'b01010 : a5 = 0;
    5'b01011 : a5 = 11;
    5'b01100 : a5 = 0;
    5'b01101 : a5 = -12;
    5'b01110 : a5 = 0;
    5'b01111 : a5 = 12;
    5'b10000 : a5 = 0;
    5'b10001 : a5 = -10;
    5'b10010 : a5 = 0;
    5'b10011 : a5 = 10;
    5'b10100 : a5 = 0;
    5'b10101 : a5 = -6;
    5'b10110 : a5 = 0;
    5'b10111 : a5 = 6;
    5'b11000 : a5 = 0;
    5'b11001 : a5 = -1;
    5'b11010 : a5 = 0;
    5'b11011 : a5 = 1;
    5'b11100 : a5 = 0;
    5'b11101 : a5 = 3;
    5'b11110 : a5 = 0;
    5'b11111 : a5 = -3;
  endcase

  a6 = 0;
  case ({STAGE[3:1], INPUT[13:12]})
    5'b00000 : a6 = 0;
    5'b00001 : a6 = -7;
    5'b00010 : a6 = 0;
    5'b00011 : a6 = 7;
    5'b00100 : a6 = 0;
    5'b00101 : a6 = -1;
    5'b00110 : a6 = 0;
    5'b00111 : a6 = 1;
    5'b01000 : a6 = 0;
    5'b01001 : a6 = 5;
    5'b01010 : a6 = 0;
    5'b01011 : a6 = -5;
    5'b01100 : a6 = 0;
    5'b01101 : a6 = 10;
    5'b01110 : a6 = 0;
    5'b01111 : a6 = -10;
    5'b10000 : a6 = 0;
    5'b10001 : a6 = 13;
    5'b10010 : a6 = 0;
    5'b10011 : a6 = -13;
    5'b10100 : a6 = 0;
    5'b10101 : a6 = 12;
    5'b10110 : a6 = 0;
    5'b10111 : a6 = -12;
    5'b11000 : a6 = 0;
    5'b11001 : a6 = 9;
    5'b11010 : a6 = 0;
    5'b11011 : a6 = -9;
    5'b11100 : a6 = 0;
    5'b11101 : a6 = 3;
    5'b11110 : a6 = 0;
    5'b11111 : a6 = -3;
  endcase

  a7 = 0;
  case ({STAGE[3:1], INPUT[15:14]})
    5'b00000 : a7 = 0;
    5'b00001 : a7 = 18;
    5'b00010 : a7 = 0;
    5'b00011 : a7 = -18;
    5'b00100 : a7 = 0;
    5'b00101 : a7 = 14;
    5'b00110 : a7 = 0;
    5'b00111 : a7 = -14;
    5'b01000 : a7 = 0;
    5'b01001 : a7 = 7;
    5'b01010 : a7 = 0;
    5'b01011 : a7 = -7;
    5'b01100 : a7 = 0;
    5'b01101 : a7 = 0;
    5'b01110 : a7 = 0;
    5'b01111 : a7 = 0;
    5'b10000 : a7 = 0;
    5'b10001 : a7 = -7;
    5'b10010 : a7 = 0;
    5'b10011 : a7 = 7;
    5'b10100 : a7 = 0;
    5'b10101 : a7 = -12;
    5'b10110 : a7 = 0;
    5'b10111 : a7 = 12;
    5'b11000 : a7 = 0;
    5'b11001 : a7 = -14;
    5'b11010 : a7 = 0;
    5'b11011 : a7 = 14;
    5'b11100 : a7 = 0;
    5'b11101 : a7 = -12;
    5'b11110 : a7 = 0;
    5'b11111 : a7 = 12;
  endcase

  a8 = 0;
  case ({STAGE[3:1], INPUT[17:16]})
    5'b00000 : a8 = 0;
    5'b00001 : a8 = -22;
    5'b00010 : a8 = 0;
    5'b00011 : a8 = 22;
    5'b00100 : a8 = 0;
    5'b00101 : a8 = -25;
    5'b00110 : a8 = 0;
    5'b00111 : a8 = 25;
    5'b01000 : a8 = 0;
    5'b01001 : a8 = -22;
    5'b01010 : a8 = 0;
    5'b01011 : a8 = 22;
    5'b01100 : a8 = 0;
    5'b01101 : a8 = -15;
    5'b01110 : a8 = 0;
    5'b01111 : a8 = 15;
    5'b10000 : a8 = 0;
    5'b10001 : a8 = -5;
    5'b10010 : a8 = 0;
    5'b10011 : a8 = 5;
    5'b10100 : a8 = 0;
    5'b10101 : a8 = 4;
    5'b10110 : a8 = 0;
    5'b10111 : a8 = -4;
    5'b11000 : a8 = 0;
    5'b11001 : a8 = 12;
    5'b11010 : a8 = 0;
    5'b11011 : a8 = -12;
    5'b11100 : a8 = 0;
    5'b11101 : a8 = 17;
    5'b11110 : a8 = 0;
    5'b11111 : a8 = -17;
  endcase

  a9 = 0;
  case ({STAGE[3:1], INPUT[19:18]})
    5'b00000 : a9 = 0;
    5'b00001 : a9 = 15;
    5'b00010 : a9 = 0;
    5'b00011 : a9 = -15;
    5'b00100 : a9 = 0;
    5'b00101 : a9 = 27;
    5'b00110 : a9 = 0;
    5'b00111 : a9 = -27;
    5'b01000 : a9 = 0;
    5'b01001 : a9 = 32;
    5'b01010 : a9 = 0;
    5'b01011 : a9 = -32;
    5'b01100 : a9 = 0;
    5'b01101 : a9 = 31;
    5'b01110 : a9 = 0;
    5'b01111 : a9 = -31;
    5'b10000 : a9 = 0;
    5'b10001 : a9 = 23;
    5'b10010 : a9 = 0;
    5'b10011 : a9 = -23;
    5'b10100 : a9 = 0;
    5'b10101 : a9 = 11;
    5'b10110 : a9 = 0;
    5'b10111 : a9 = -11;
    5'b11000 : a9 = 0;
    5'b11001 : a9 = -2;
    5'b11010 : a9 = 0;
    5'b11011 : a9 = 2;
    5'b11100 : a9 = 0;
    5'b11101 : a9 = -14;
    5'b11110 : a9 = 0;
    5'b11111 : a9 = 14;
  endcase

  a10 = 0;
  case ({STAGE[3:1], INPUT[21:20]})
    5'b00000 : a10 = 0;
    5'b00001 : a10 = 8;
    5'b00010 : a10 = 0;
    5'b00011 : a10 = -8;
    5'b00100 : a10 = 0;
    5'b00101 : a10 = -10;
    5'b00110 : a10 = 0;
    5'b00111 : a10 = 10;
    5'b01000 : a10 = 0;
    5'b01001 : a10 = -26;
    5'b01010 : a10 = 0;
    5'b01011 : a10 = 26;
    5'b01100 : a10 = 0;
    5'b01101 : a10 = -35;
    5'b01110 : a10 = 0;
    5'b01111 : a10 = 35;
    5'b10000 : a10 = 0;
    5'b10001 : a10 = -36;
    5'b10010 : a10 = 0;
    5'b10011 : a10 = 36;
    5'b10100 : a10 = 0;
    5'b10101 : a10 = -29;
    5'b10110 : a10 = 0;
    5'b10111 : a10 = 29;
    5'b11000 : a10 = 0;
    5'b11001 : a10 = -16;
    5'b11010 : a10 = 0;
    5'b11011 : a10 = 16;
    5'b11100 : a10 = 0;
    5'b11101 : a10 = 0;
    5'b11110 : a10 = 0;
    5'b11111 : a10 = 0;
  endcase

  a11 = 0;
  case ({STAGE[3:1], INPUT[23:22]})
    5'b00000 : a11 = 0;
    5'b00001 : a11 = -50;
    5'b00010 : a11 = 0;
    5'b00011 : a11 = 50;
    5'b00100 : a11 = 0;
    5'b00101 : a11 = -32;
    5'b00110 : a11 = 0;
    5'b00111 : a11 = 32;
    5'b01000 : a11 = 0;
    5'b01001 : a11 = -9;
    5'b01010 : a11 = 0;
    5'b01011 : a11 = 9;
    5'b01100 : a11 = 0;
    5'b01101 : a11 = 14;
    5'b01110 : a11 = 0;
    5'b01111 : a11 = -14;
    5'b10000 : a11 = 0;
    5'b10001 : a11 = 31;
    5'b10010 : a11 = 0;
    5'b10011 : a11 = -31;
    5'b10100 : a11 = 0;
    5'b10101 : a11 = 39;
    5'b10110 : a11 = 0;
    5'b10111 : a11 = -39;
    5'b11000 : a11 = 0;
    5'b11001 : a11 = 37;
    5'b11010 : a11 = 0;
    5'b11011 : a11 = -37;
    5'b11100 : a11 = 0;
    5'b11101 : a11 = 26;
    5'b11110 : a11 = 0;
    5'b11111 : a11 = -26;
  endcase

  a12 = 0;
  case ({STAGE[3:1], INPUT[25:24]})
    5'b00000 : a12 = 0;
    5'b00001 : a12 = 105;
    5'b00010 : a12 = 0;
    5'b00011 : a12 = -105;
    5'b00100 : a12 = 0;
    5'b00101 : a12 = 106;
    5'b00110 : a12 = 0;
    5'b00111 : a12 = -106;
    5'b01000 : a12 = 0;
    5'b01001 : a12 = 85;
    5'b01010 : a12 = 0;
    5'b01011 : a12 = -85;
    5'b01100 : a12 = 0;
    5'b01101 : a12 = 49;
    5'b01110 : a12 = 0;
    5'b01111 : a12 = -49;
    5'b10000 : a12 = 0;
    5'b10001 : a12 = 10;
    5'b10010 : a12 = 0;
    5'b10011 : a12 = -10;
    5'b10100 : a12 = 0;
    5'b10101 : a12 = -24;
    5'b10110 : a12 = 0;
    5'b10111 : a12 = 24;
    5'b11000 : a12 = 0;
    5'b11001 : a12 = -48;
    5'b11010 : a12 = 0;
    5'b11011 : a12 = 48;
    5'b11100 : a12 = 0;
    5'b11101 : a12 = -56;
    5'b11110 : a12 = 0;
    5'b11111 : a12 = 56;
  endcase

  a13 = 0;
  case ({STAGE[3:1], INPUT[27:26]})
    5'b00000 : a13 = 0;
    5'b00001 : a13 = -166;
    5'b00010 : a13 = 0;
    5'b00011 : a13 = 166;
    5'b00100 : a13 = 0;
    5'b00101 : a13 = -214;
    5'b00110 : a13 = 0;
    5'b00111 : a13 = 214;
    5'b01000 : a13 = 0;
    5'b01001 : a13 = -215;
    5'b01010 : a13 = 0;
    5'b01011 : a13 = 215;
    5'b01100 : a13 = 0;
    5'b01101 : a13 = -177;
    5'b01110 : a13 = 0;
    5'b01111 : a13 = 177;
    5'b10000 : a13 = 0;
    5'b10001 : a13 = -113;
    5'b10010 : a13 = 0;
    5'b10011 : a13 = 113;
    5'b10100 : a13 = 0;
    5'b10101 : a13 = -39;
    5'b10110 : a13 = 0;
    5'b10111 : a13 = 39;
    5'b11000 : a13 = 0;
    5'b11001 : a13 = 28;
    5'b11010 : a13 = 0;
    5'b11011 : a13 = -28;
    5'b11100 : a13 = 0;
    5'b11101 : a13 = 79;
    5'b11110 : a13 = 0;
    5'b11111 : a13 = -79;
  endcase

  a14 = 0;
  case ({STAGE[3:1], INPUT[29:28]})
    5'b00000 : a14 = 0;
    5'b00001 : a14 = 222;
    5'b00010 : a14 = 0;
    5'b00011 : a14 = -222;
    5'b00100 : a14 = 0;
    5'b00101 : a14 = 370;
    5'b00110 : a14 = 0;
    5'b00111 : a14 = -370;
    5'b01000 : a14 = 0;
    5'b01001 : a14 = 431;
    5'b01010 : a14 = 0;
    5'b01011 : a14 = -431;
    5'b01100 : a14 = 0;
    5'b01101 : a14 = 408;
    5'b01110 : a14 = 0;
    5'b01111 : a14 = -408;
    5'b10000 : a14 = 0;
    5'b10001 : a14 = 320;
    5'b10010 : a14 = 0;
    5'b10011 : a14 = -320;
    5'b10100 : a14 = 0;
    5'b10101 : a14 = 192;
    5'b10110 : a14 = 0;
    5'b10111 : a14 = -192;
    5'b11000 : a14 = 0;
    5'b11001 : a14 = 51;
    5'b11010 : a14 = 0;
    5'b11011 : a14 = -51;
    5'b11100 : a14 = 0;
    5'b11101 : a14 = -74;
    5'b11110 : a14 = 0;
    5'b11111 : a14 = 74;
  endcase

  a15 = 0;
  case ({STAGE[3:1], INPUT[31:30]})
    5'b00000 : a15 = 0;
    5'b00001 : a15 = -261;
    5'b00010 : a15 = 0;
    5'b00011 : a15 = 261;
    5'b00100 : a15 = 0;
    5'b00101 : a15 = -665;
    5'b00110 : a15 = 0;
    5'b00111 : a15 = 665;
    5'b01000 : a15 = 0;
    5'b01001 : a15 = -873;
    5'b01010 : a15 = 0;
    5'b01011 : a15 = 873;
    5'b01100 : a15 = 0;
    5'b01101 : a15 = -897;
    5'b01110 : a15 = 0;
    5'b01111 : a15 = 897;
    5'b10000 : a15 = 0;
    5'b10001 : a15 = -771;
    5'b10010 : a15 = 0;
    5'b10011 : a15 = 771;
    5'b10100 : a15 = 0;
    5'b10101 : a15 = -545;
    5'b10110 : a15 = 0;
    5'b10111 : a15 = 545;
    5'b11000 : a15 = 0;
    5'b11001 : a15 = -270;
    5'b11010 : a15 = 0;
    5'b11011 : a15 = 270;
    5'b11100 : a15 = 0;
    5'b11101 : a15 = 0;
    5'b11110 : a15 = 0;
    5'b11111 : a15 = 0;
  endcase

  a16 = 0;
  case ({STAGE[3:1], INPUT[33:32]})
    5'b00000 : a16 = 0;
    5'b00001 : a16 = 4651;
    5'b00010 : a16 = 0;
    5'b00011 : a16 = -4651;
    5'b00100 : a16 = 0;
    5'b00101 : a16 = 4513;
    5'b00110 : a16 = 0;
    5'b00111 : a16 = -4513;
    5'b01000 : a16 = 0;
    5'b01001 : a16 = 4114;
    5'b01010 : a16 = 0;
    5'b01011 : a16 = -4114;
    5'b01100 : a16 = 0;
    5'b01101 : a16 = 3498;
    5'b01110 : a16 = 0;
    5'b01111 : a16 = -3498;
    5'b10000 : a16 = 0;
    5'b10001 : a16 = 2731;
    5'b10010 : a16 = 0;
    5'b10011 : a16 = -2731;
    5'b10100 : a16 = 0;
    5'b10101 : a16 = 1892;
    5'b10110 : a16 = 0;
    5'b10111 : a16 = -1892;
    5'b11000 : a16 = 0;
    5'b11001 : a16 = 1066;
    5'b11010 : a16 = 0;
    5'b11011 : a16 = -1066;
    5'b11100 : a16 = 0;
    5'b11101 : a16 = 328;
    5'b11110 : a16 = 0;
    5'b11111 : a16 = -328;
  endcase

  a17 = 0;
  case ({STAGE[3:1], INPUT[35:34]})
    5'b00000 : a17 = 0;
    5'b00001 : a17 = -261;
    5'b00010 : a17 = 0;
    5'b00011 : a17 = 261;
    5'b00100 : a17 = 0;
    5'b00101 : a17 = 328;
    5'b00110 : a17 = 0;
    5'b00111 : a17 = -328;
    5'b01000 : a17 = 0;
    5'b01001 : a17 = 1066;
    5'b01010 : a17 = 0;
    5'b01011 : a17 = -1066;
    5'b01100 : a17 = 0;
    5'b01101 : a17 = 1892;
    5'b01110 : a17 = 0;
    5'b01111 : a17 = -1892;
    5'b10000 : a17 = 0;
    5'b10001 : a17 = 2731;
    5'b10010 : a17 = 0;
    5'b10011 : a17 = -2731;
    5'b10100 : a17 = 0;
    5'b10101 : a17 = 3498;
    5'b10110 : a17 = 0;
    5'b10111 : a17 = -3498;
    5'b11000 : a17 = 0;
    5'b11001 : a17 = 4114;
    5'b11010 : a17 = 0;
    5'b11011 : a17 = -4114;
    5'b11100 : a17 = 0;
    5'b11101 : a17 = 4513;
    5'b11110 : a17 = 0;
    5'b11111 : a17 = -4513;
  endcase

  a18 = 0;
  case ({STAGE[3:1], INPUT[37:36]})
    5'b00000 : a18 = 0;
    5'b00001 : a18 = 222;
    5'b00010 : a18 = 0;
    5'b00011 : a18 = -222;
    5'b00100 : a18 = 0;
    5'b00101 : a18 = 0;
    5'b00110 : a18 = 0;
    5'b00111 : a18 = 0;
    5'b01000 : a18 = 0;
    5'b01001 : a18 = -270;
    5'b01010 : a18 = 0;
    5'b01011 : a18 = 270;
    5'b01100 : a18 = 0;
    5'b01101 : a18 = -545;
    5'b01110 : a18 = 0;
    5'b01111 : a18 = 545;
    5'b10000 : a18 = 0;
    5'b10001 : a18 = -771;
    5'b10010 : a18 = 0;
    5'b10011 : a18 = 771;
    5'b10100 : a18 = 0;
    5'b10101 : a18 = -897;
    5'b10110 : a18 = 0;
    5'b10111 : a18 = 897;
    5'b11000 : a18 = 0;
    5'b11001 : a18 = -873;
    5'b11010 : a18 = 0;
    5'b11011 : a18 = 873;
    5'b11100 : a18 = 0;
    5'b11101 : a18 = -665;
    5'b11110 : a18 = 0;
    5'b11111 : a18 = 665;
  endcase

  a19 = 0;
  case ({STAGE[3:1], INPUT[39:38]})
    5'b00000 : a19 = 0;
    5'b00001 : a19 = -166;
    5'b00010 : a19 = 0;
    5'b00011 : a19 = 166;
    5'b00100 : a19 = 0;
    5'b00101 : a19 = -74;
    5'b00110 : a19 = 0;
    5'b00111 : a19 = 74;
    5'b01000 : a19 = 0;
    5'b01001 : a19 = 51;
    5'b01010 : a19 = 0;
    5'b01011 : a19 = -51;
    5'b01100 : a19 = 0;
    5'b01101 : a19 = 192;
    5'b01110 : a19 = 0;
    5'b01111 : a19 = -192;
    5'b10000 : a19 = 0;
    5'b10001 : a19 = 320;
    5'b10010 : a19 = 0;
    5'b10011 : a19 = -320;
    5'b10100 : a19 = 0;
    5'b10101 : a19 = 408;
    5'b10110 : a19 = 0;
    5'b10111 : a19 = -408;
    5'b11000 : a19 = 0;
    5'b11001 : a19 = 431;
    5'b11010 : a19 = 0;
    5'b11011 : a19 = -431;
    5'b11100 : a19 = 0;
    5'b11101 : a19 = 370;
    5'b11110 : a19 = 0;
    5'b11111 : a19 = -370;
  endcase

  a20 = 0;
  case ({STAGE[3:1], INPUT[41:40]})
    5'b00000 : a20 = 0;
    5'b00001 : a20 = 105;
    5'b00010 : a20 = 0;
    5'b00011 : a20 = -105;
    5'b00100 : a20 = 0;
    5'b00101 : a20 = 79;
    5'b00110 : a20 = 0;
    5'b00111 : a20 = -79;
    5'b01000 : a20 = 0;
    5'b01001 : a20 = 28;
    5'b01010 : a20 = 0;
    5'b01011 : a20 = -28;
    5'b01100 : a20 = 0;
    5'b01101 : a20 = -39;
    5'b01110 : a20 = 0;
    5'b01111 : a20 = 39;
    5'b10000 : a20 = 0;
    5'b10001 : a20 = -113;
    5'b10010 : a20 = 0;
    5'b10011 : a20 = 113;
    5'b10100 : a20 = 0;
    5'b10101 : a20 = -177;
    5'b10110 : a20 = 0;
    5'b10111 : a20 = 177;
    5'b11000 : a20 = 0;
    5'b11001 : a20 = -215;
    5'b11010 : a20 = 0;
    5'b11011 : a20 = 215;
    5'b11100 : a20 = 0;
    5'b11101 : a20 = -214;
    5'b11110 : a20 = 0;
    5'b11111 : a20 = 214;
  endcase

  a21 = 0;
  case ({STAGE[3:1], INPUT[43:42]})
    5'b00000 : a21 = 0;
    5'b00001 : a21 = -50;
    5'b00010 : a21 = 0;
    5'b00011 : a21 = 50;
    5'b00100 : a21 = 0;
    5'b00101 : a21 = -56;
    5'b00110 : a21 = 0;
    5'b00111 : a21 = 56;
    5'b01000 : a21 = 0;
    5'b01001 : a21 = -48;
    5'b01010 : a21 = 0;
    5'b01011 : a21 = 48;
    5'b01100 : a21 = 0;
    5'b01101 : a21 = -24;
    5'b01110 : a21 = 0;
    5'b01111 : a21 = 24;
    5'b10000 : a21 = 0;
    5'b10001 : a21 = 10;
    5'b10010 : a21 = 0;
    5'b10011 : a21 = -10;
    5'b10100 : a21 = 0;
    5'b10101 : a21 = 49;
    5'b10110 : a21 = 0;
    5'b10111 : a21 = -49;
    5'b11000 : a21 = 0;
    5'b11001 : a21 = 85;
    5'b11010 : a21 = 0;
    5'b11011 : a21 = -85;
    5'b11100 : a21 = 0;
    5'b11101 : a21 = 106;
    5'b11110 : a21 = 0;
    5'b11111 : a21 = -106;
  endcase

  a22 = 0;
  case ({STAGE[3:1], INPUT[45:44]})
    5'b00000 : a22 = 0;
    5'b00001 : a22 = 8;
    5'b00010 : a22 = 0;
    5'b00011 : a22 = -8;
    5'b00100 : a22 = 0;
    5'b00101 : a22 = 26;
    5'b00110 : a22 = 0;
    5'b00111 : a22 = -26;
    5'b01000 : a22 = 0;
    5'b01001 : a22 = 37;
    5'b01010 : a22 = 0;
    5'b01011 : a22 = -37;
    5'b01100 : a22 = 0;
    5'b01101 : a22 = 39;
    5'b01110 : a22 = 0;
    5'b01111 : a22 = -39;
    5'b10000 : a22 = 0;
    5'b10001 : a22 = 31;
    5'b10010 : a22 = 0;
    5'b10011 : a22 = -31;
    5'b10100 : a22 = 0;
    5'b10101 : a22 = 14;
    5'b10110 : a22 = 0;
    5'b10111 : a22 = -14;
    5'b11000 : a22 = 0;
    5'b11001 : a22 = -9;
    5'b11010 : a22 = 0;
    5'b11011 : a22 = 9;
    5'b11100 : a22 = 0;
    5'b11101 : a22 = -32;
    5'b11110 : a22 = 0;
    5'b11111 : a22 = 32;
  endcase

  a23 = 0;
  case ({STAGE[3:1], INPUT[47:46]})
    5'b00000 : a23 = 0;
    5'b00001 : a23 = 15;
    5'b00010 : a23 = 0;
    5'b00011 : a23 = -15;
    5'b00100 : a23 = 0;
    5'b00101 : a23 = 0;
    5'b00110 : a23 = 0;
    5'b00111 : a23 = 0;
    5'b01000 : a23 = 0;
    5'b01001 : a23 = -16;
    5'b01010 : a23 = 0;
    5'b01011 : a23 = 16;
    5'b01100 : a23 = 0;
    5'b01101 : a23 = -29;
    5'b01110 : a23 = 0;
    5'b01111 : a23 = 29;
    5'b10000 : a23 = 0;
    5'b10001 : a23 = -36;
    5'b10010 : a23 = 0;
    5'b10011 : a23 = 36;
    5'b10100 : a23 = 0;
    5'b10101 : a23 = -35;
    5'b10110 : a23 = 0;
    5'b10111 : a23 = 35;
    5'b11000 : a23 = 0;
    5'b11001 : a23 = -26;
    5'b11010 : a23 = 0;
    5'b11011 : a23 = 26;
    5'b11100 : a23 = 0;
    5'b11101 : a23 = -10;
    5'b11110 : a23 = 0;
    5'b11111 : a23 = 10;
  endcase

  a24 = 0;
  case ({STAGE[3:1], INPUT[49:48]})
    5'b00000 : a24 = 0;
    5'b00001 : a24 = -22;
    5'b00010 : a24 = 0;
    5'b00011 : a24 = 22;
    5'b00100 : a24 = 0;
    5'b00101 : a24 = -14;
    5'b00110 : a24 = 0;
    5'b00111 : a24 = 14;
    5'b01000 : a24 = 0;
    5'b01001 : a24 = -2;
    5'b01010 : a24 = 0;
    5'b01011 : a24 = 2;
    5'b01100 : a24 = 0;
    5'b01101 : a24 = 11;
    5'b01110 : a24 = 0;
    5'b01111 : a24 = -11;
    5'b10000 : a24 = 0;
    5'b10001 : a24 = 23;
    5'b10010 : a24 = 0;
    5'b10011 : a24 = -23;
    5'b10100 : a24 = 0;
    5'b10101 : a24 = 31;
    5'b10110 : a24 = 0;
    5'b10111 : a24 = -31;
    5'b11000 : a24 = 0;
    5'b11001 : a24 = 32;
    5'b11010 : a24 = 0;
    5'b11011 : a24 = -32;
    5'b11100 : a24 = 0;
    5'b11101 : a24 = 27;
    5'b11110 : a24 = 0;
    5'b11111 : a24 = -27;
  endcase

  a25 = 0;
  case ({STAGE[3:1], INPUT[51:50]})
    5'b00000 : a25 = 0;
    5'b00001 : a25 = 18;
    5'b00010 : a25 = 0;
    5'b00011 : a25 = -18;
    5'b00100 : a25 = 0;
    5'b00101 : a25 = 17;
    5'b00110 : a25 = 0;
    5'b00111 : a25 = -17;
    5'b01000 : a25 = 0;
    5'b01001 : a25 = 12;
    5'b01010 : a25 = 0;
    5'b01011 : a25 = -12;
    5'b01100 : a25 = 0;
    5'b01101 : a25 = 4;
    5'b01110 : a25 = 0;
    5'b01111 : a25 = -4;
    5'b10000 : a25 = 0;
    5'b10001 : a25 = -5;
    5'b10010 : a25 = 0;
    5'b10011 : a25 = 5;
    5'b10100 : a25 = 0;
    5'b10101 : a25 = -15;
    5'b10110 : a25 = 0;
    5'b10111 : a25 = 15;
    5'b11000 : a25 = 0;
    5'b11001 : a25 = -22;
    5'b11010 : a25 = 0;
    5'b11011 : a25 = 22;
    5'b11100 : a25 = 0;
    5'b11101 : a25 = -25;
    5'b11110 : a25 = 0;
    5'b11111 : a25 = 25;
  endcase

  a26 = 0;
  case ({STAGE[3:1], INPUT[53:52]})
    5'b00000 : a26 = 0;
    5'b00001 : a26 = -7;
    5'b00010 : a26 = 0;
    5'b00011 : a26 = 7;
    5'b00100 : a26 = 0;
    5'b00101 : a26 = -12;
    5'b00110 : a26 = 0;
    5'b00111 : a26 = 12;
    5'b01000 : a26 = 0;
    5'b01001 : a26 = -14;
    5'b01010 : a26 = 0;
    5'b01011 : a26 = 14;
    5'b01100 : a26 = 0;
    5'b01101 : a26 = -12;
    5'b01110 : a26 = 0;
    5'b01111 : a26 = 12;
    5'b10000 : a26 = 0;
    5'b10001 : a26 = -7;
    5'b10010 : a26 = 0;
    5'b10011 : a26 = 7;
    5'b10100 : a26 = 0;
    5'b10101 : a26 = 0;
    5'b10110 : a26 = 0;
    5'b10111 : a26 = 0;
    5'b11000 : a26 = 0;
    5'b11001 : a26 = 7;
    5'b11010 : a26 = 0;
    5'b11011 : a26 = -7;
    5'b11100 : a26 = 0;
    5'b11101 : a26 = 14;
    5'b11110 : a26 = 0;
    5'b11111 : a26 = -14;
  endcase

  a27 = 0;
  case ({STAGE[3:1], INPUT[55:54]})
    5'b00000 : a27 = 0;
    5'b00001 : a27 = -2;
    5'b00010 : a27 = 0;
    5'b00011 : a27 = 2;
    5'b00100 : a27 = 0;
    5'b00101 : a27 = 3;
    5'b00110 : a27 = 0;
    5'b00111 : a27 = -3;
    5'b01000 : a27 = 0;
    5'b01001 : a27 = 9;
    5'b01010 : a27 = 0;
    5'b01011 : a27 = -9;
    5'b01100 : a27 = 0;
    5'b01101 : a27 = 12;
    5'b01110 : a27 = 0;
    5'b01111 : a27 = -12;
    5'b10000 : a27 = 0;
    5'b10001 : a27 = 13;
    5'b10010 : a27 = 0;
    5'b10011 : a27 = -13;
    5'b10100 : a27 = 0;
    5'b10101 : a27 = 10;
    5'b10110 : a27 = 0;
    5'b10111 : a27 = -10;
    5'b11000 : a27 = 0;
    5'b11001 : a27 = 5;
    5'b11010 : a27 = 0;
    5'b11011 : a27 = -5;
    5'b11100 : a27 = 0;
    5'b11101 : a27 = -1;
    5'b11110 : a27 = 0;
    5'b11111 : a27 = 1;
  endcase

  a28 = 0;
  case ({STAGE[3:1], INPUT[57:56]})
    5'b00000 : a28 = 0;
    5'b00001 : a28 = 8;
    5'b00010 : a28 = 0;
    5'b00011 : a28 = -8;
    5'b00100 : a28 = 0;
    5'b00101 : a28 = 3;
    5'b00110 : a28 = 0;
    5'b00111 : a28 = -3;
    5'b01000 : a28 = 0;
    5'b01001 : a28 = -1;
    5'b01010 : a28 = 0;
    5'b01011 : a28 = 1;
    5'b01100 : a28 = 0;
    5'b01101 : a28 = -6;
    5'b01110 : a28 = 0;
    5'b01111 : a28 = 6;
    5'b10000 : a28 = 0;
    5'b10001 : a28 = -10;
    5'b10010 : a28 = 0;
    5'b10011 : a28 = 10;
    5'b10100 : a28 = 0;
    5'b10101 : a28 = -12;
    5'b10110 : a28 = 0;
    5'b10111 : a28 = 12;
    5'b11000 : a28 = 0;
    5'b11001 : a28 = -11;
    5'b11010 : a28 = 0;
    5'b11011 : a28 = 11;
    5'b11100 : a28 = 0;
    5'b11101 : a28 = -7;
    5'b11110 : a28 = 0;
    5'b11111 : a28 = 7;
  endcase

  a29 = 0;
  case ({STAGE[3:1], INPUT[59:58]})
    5'b00000 : a29 = 0;
    5'b00001 : a29 = -9;
    5'b00010 : a29 = 0;
    5'b00011 : a29 = 9;
    5'b00100 : a29 = 0;
    5'b00101 : a29 = -7;
    5'b00110 : a29 = 0;
    5'b00111 : a29 = 7;
    5'b01000 : a29 = 0;
    5'b01001 : a29 = -4;
    5'b01010 : a29 = 0;
    5'b01011 : a29 = 4;
    5'b01100 : a29 = 0;
    5'b01101 : a29 = 0;
    5'b01110 : a29 = 0;
    5'b01111 : a29 = 0;
    5'b10000 : a29 = 0;
    5'b10001 : a29 = 4;
    5'b10010 : a29 = 0;
    5'b10011 : a29 = -4;
    5'b10100 : a29 = 0;
    5'b10101 : a29 = 8;
    5'b10110 : a29 = 0;
    5'b10111 : a29 = -8;
    5'b11000 : a29 = 0;
    5'b11001 : a29 = 10;
    5'b11010 : a29 = 0;
    5'b11011 : a29 = -10;
    5'b11100 : a29 = 0;
    5'b11101 : a29 = 10;
    5'b11110 : a29 = 0;
    5'b11111 : a29 = -10;
  endcase

  a30 = 0;
  case ({STAGE[3:1], INPUT[61:60]})
    5'b00000 : a30 = 0;
    5'b00001 : a30 = 5;
    5'b00010 : a30 = 0;
    5'b00011 : a30 = -5;
    5'b00100 : a30 = 0;
    5'b00101 : a30 = 7;
    5'b00110 : a30 = 0;
    5'b00111 : a30 = -7;
    5'b01000 : a30 = 0;
    5'b01001 : a30 = 7;
    5'b01010 : a30 = 0;
    5'b01011 : a30 = -7;
    5'b01100 : a30 = 0;
    5'b01101 : a30 = 5;
    5'b01110 : a30 = 0;
    5'b01111 : a30 = -5;
    5'b10000 : a30 = 0;
    5'b10001 : a30 = 2;
    5'b10010 : a30 = 0;
    5'b10011 : a30 = -2;
    5'b10100 : a30 = 0;
    5'b10101 : a30 = -1;
    5'b10110 : a30 = 0;
    5'b10111 : a30 = 1;
    5'b11000 : a30 = 0;
    5'b11001 : a30 = -5;
    5'b11010 : a30 = 0;
    5'b11011 : a30 = 5;
    5'b11100 : a30 = 0;
    5'b11101 : a30 = -8;
    5'b11110 : a30 = 0;
    5'b11111 : a30 = 8;
  endcase

  a31 = 0;
  case ({STAGE[3:1], INPUT[63:62]})
    5'b00000 : a31 = 0;
    5'b00001 : a31 = 0;
    5'b00010 : a31 = 0;
    5'b00011 : a31 = 0;
    5'b00100 : a31 = 0;
    5'b00101 : a31 = -3;
    5'b00110 : a31 = 0;
    5'b00111 : a31 = 3;
    5'b01000 : a31 = 0;
    5'b01001 : a31 = -5;
    5'b01010 : a31 = 0;
    5'b01011 : a31 = 5;
    5'b01100 : a31 = 0;
    5'b01101 : a31 = -6;
    5'b01110 : a31 = 0;
    5'b01111 : a31 = 6;
    5'b10000 : a31 = 0;
    5'b10001 : a31 = -6;
    5'b10010 : a31 = 0;
    5'b10011 : a31 = 6;
    5'b10100 : a31 = 0;
    5'b10101 : a31 = -3;
    5'b10110 : a31 = 0;
    5'b10111 : a31 = 3;
    5'b11000 : a31 = 0;
    5'b11001 : a31 = 0;
    5'b11010 : a31 = 0;
    5'b11011 : a31 = 0;
    5'b11100 : a31 = 0;
    5'b11101 : a31 = 2;
    5'b11110 : a31 = 0;
    5'b11111 : a31 = -2;
  endcase

  a32 = 0;
  case ({STAGE[3:1], INPUT[65:64]})
    5'b00000 : a32 = 0;
    5'b00001 : a32 = -3;
    5'b00010 : a32 = 0;
    5'b00011 : a32 = 3;
    5'b00100 : a32 = 0;
    5'b00101 : a32 = 0;
    5'b00110 : a32 = 0;
    5'b00111 : a32 = 0;
    5'b01000 : a32 = 0;
    5'b01001 : a32 = 2;
    5'b01010 : a32 = 0;
    5'b01011 : a32 = -2;
    5'b01100 : a32 = 0;
    5'b01101 : a32 = 4;
    5'b01110 : a32 = 0;
    5'b01111 : a32 = -4;
    5'b10000 : a32 = 0;
    5'b10001 : a32 = 6;
    5'b10010 : a32 = 0;
    5'b10011 : a32 = -6;
    5'b10100 : a32 = 0;
    5'b10101 : a32 = 6;
    5'b10110 : a32 = 0;
    5'b10111 : a32 = -6;
    5'b11000 : a32 = 0;
    5'b11001 : a32 = 5;
    5'b11010 : a32 = 0;
    5'b11011 : a32 = -5;
    5'b11100 : a32 = 0;
    5'b11101 : a32 = 2;
    5'b11110 : a32 = 0;
    5'b11111 : a32 = -2;
  endcase

end
assign sum =  a0  + a1  + a2  + a3  + a4  + a5  + a6  + a7  + 
              a8  + a9  + a10 + a11 + a12 + a13 + a14 + a15 +
              a16 + a17 + a18 + a19 + a20 + a21 + a22 + a23 +
              a24 + a25 + a26 + a27 + a28 + a29 + a30 + a31 + 
              a32;

always @(posedge CLK)
  begin
    if (STAGE[0] == 0 && ENABLE)
    begin
      result_i <= sum[13:1];
      //$monitor ("%t Display OUTPUT_I : %h", $time, result_i);
    end
    else if (STAGE[0] == 1 && ENABLE)
    begin
      result_q <= sum[13:1];
     // $monitor ("%t Display OUTPUT_Q : %h", $time, result_q);
    end
  end

endmodule